* NGSPICE file created from (UNNAMED).ext - technology: minimum

.subckt UNNAMED)
.ends

